** Profile: "SCHEMATIC1-bias"  [ C:\Users\emiba\OneDrive\Desktop\P1_B_N1\proiect-sim-pspicefiles\schematic1\bias.sim ] 

** Creating circuit file "bias.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../lib_modelepspice_anexa_1_a/modele_a1_lib/bc856b.lib" 
.LIB "../../../lib_modelepspice_anexa_1_a/modele_a1_lib/bc846b.lib" 
.LIB "../../../proiect-sim-pspicefiles/schematic1/test/1n4148.lib" 
* From [PSPICE NETLIST] section of C:\Users\emiba\AppData\Roaming\SPB_16.6\cdssetup\OrCAD_PSpice\24.1.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 10ms 0 1u 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\SCHEMATIC1.net" 


.END
